module test_comm;
    initial begin
        #10;
    end
endmodule
